`timescale 1ns / 1ps

// Engineer: Tanay Das

module not_gate(
    input a,
    output b
    );
    
    assign b = ~a;
endmodule


